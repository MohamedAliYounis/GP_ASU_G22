magic
tech sky130A
magscale 1 2
timestamp 1654633061
<< obsli1 >>
rect 1104 2159 398820 397681
<< obsm1 >>
rect 1104 1368 398820 397712
<< metal2 >>
rect 3790 399200 3846 400000
rect 11426 399200 11482 400000
rect 19154 399200 19210 400000
rect 26790 399200 26846 400000
rect 34518 399200 34574 400000
rect 42246 399200 42302 400000
rect 49882 399200 49938 400000
rect 57610 399200 57666 400000
rect 65246 399200 65302 400000
rect 72974 399200 73030 400000
rect 80702 399200 80758 400000
rect 88338 399200 88394 400000
rect 96066 399200 96122 400000
rect 103794 399200 103850 400000
rect 111430 399200 111486 400000
rect 119158 399200 119214 400000
rect 126794 399200 126850 400000
rect 134522 399200 134578 400000
rect 142250 399200 142306 400000
rect 149886 399200 149942 400000
rect 157614 399200 157670 400000
rect 165250 399200 165306 400000
rect 172978 399200 173034 400000
rect 180706 399200 180762 400000
rect 188342 399200 188398 400000
rect 196070 399200 196126 400000
rect 203798 399200 203854 400000
rect 211434 399200 211490 400000
rect 219162 399200 219218 400000
rect 226798 399200 226854 400000
rect 234526 399200 234582 400000
rect 242254 399200 242310 400000
rect 249890 399200 249946 400000
rect 257618 399200 257674 400000
rect 265254 399200 265310 400000
rect 272982 399200 273038 400000
rect 280710 399200 280766 400000
rect 288346 399200 288402 400000
rect 296074 399200 296130 400000
rect 303802 399200 303858 400000
rect 311438 399200 311494 400000
rect 319166 399200 319222 400000
rect 326802 399200 326858 400000
rect 334530 399200 334586 400000
rect 342258 399200 342314 400000
rect 349894 399200 349950 400000
rect 357622 399200 357678 400000
rect 365258 399200 365314 400000
rect 372986 399200 373042 400000
rect 380714 399200 380770 400000
rect 388350 399200 388406 400000
rect 396078 399200 396134 400000
rect 2778 0 2834 800
rect 8390 0 8446 800
rect 14002 0 14058 800
rect 19614 0 19670 800
rect 25226 0 25282 800
rect 30930 0 30986 800
rect 36542 0 36598 800
rect 42154 0 42210 800
rect 47766 0 47822 800
rect 53470 0 53526 800
rect 59082 0 59138 800
rect 64694 0 64750 800
rect 70306 0 70362 800
rect 76010 0 76066 800
rect 81622 0 81678 800
rect 87234 0 87290 800
rect 92846 0 92902 800
rect 98550 0 98606 800
rect 104162 0 104218 800
rect 109774 0 109830 800
rect 115386 0 115442 800
rect 121090 0 121146 800
rect 126702 0 126758 800
rect 132314 0 132370 800
rect 137926 0 137982 800
rect 143538 0 143594 800
rect 149242 0 149298 800
rect 154854 0 154910 800
rect 160466 0 160522 800
rect 166078 0 166134 800
rect 171782 0 171838 800
rect 177394 0 177450 800
rect 183006 0 183062 800
rect 188618 0 188674 800
rect 194322 0 194378 800
rect 199934 0 199990 800
rect 205546 0 205602 800
rect 211158 0 211214 800
rect 216862 0 216918 800
rect 222474 0 222530 800
rect 228086 0 228142 800
rect 233698 0 233754 800
rect 239402 0 239458 800
rect 245014 0 245070 800
rect 250626 0 250682 800
rect 256238 0 256294 800
rect 261942 0 261998 800
rect 267554 0 267610 800
rect 273166 0 273222 800
rect 278778 0 278834 800
rect 284390 0 284446 800
rect 290094 0 290150 800
rect 295706 0 295762 800
rect 301318 0 301374 800
rect 306930 0 306986 800
rect 312634 0 312690 800
rect 318246 0 318302 800
rect 323858 0 323914 800
rect 329470 0 329526 800
rect 335174 0 335230 800
rect 340786 0 340842 800
rect 346398 0 346454 800
rect 352010 0 352066 800
rect 357714 0 357770 800
rect 363326 0 363382 800
rect 368938 0 368994 800
rect 374550 0 374606 800
rect 380254 0 380310 800
rect 385866 0 385922 800
rect 391478 0 391534 800
rect 397090 0 397146 800
<< obsm2 >>
rect 1398 399144 3734 399242
rect 3902 399144 11370 399242
rect 11538 399144 19098 399242
rect 19266 399144 26734 399242
rect 26902 399144 34462 399242
rect 34630 399144 42190 399242
rect 42358 399144 49826 399242
rect 49994 399144 57554 399242
rect 57722 399144 65190 399242
rect 65358 399144 72918 399242
rect 73086 399144 80646 399242
rect 80814 399144 88282 399242
rect 88450 399144 96010 399242
rect 96178 399144 103738 399242
rect 103906 399144 111374 399242
rect 111542 399144 119102 399242
rect 119270 399144 126738 399242
rect 126906 399144 134466 399242
rect 134634 399144 142194 399242
rect 142362 399144 149830 399242
rect 149998 399144 157558 399242
rect 157726 399144 165194 399242
rect 165362 399144 172922 399242
rect 173090 399144 180650 399242
rect 180818 399144 188286 399242
rect 188454 399144 196014 399242
rect 196182 399144 203742 399242
rect 203910 399144 211378 399242
rect 211546 399144 219106 399242
rect 219274 399144 226742 399242
rect 226910 399144 234470 399242
rect 234638 399144 242198 399242
rect 242366 399144 249834 399242
rect 250002 399144 257562 399242
rect 257730 399144 265198 399242
rect 265366 399144 272926 399242
rect 273094 399144 280654 399242
rect 280822 399144 288290 399242
rect 288458 399144 296018 399242
rect 296186 399144 303746 399242
rect 303914 399144 311382 399242
rect 311550 399144 319110 399242
rect 319278 399144 326746 399242
rect 326914 399144 334474 399242
rect 334642 399144 342202 399242
rect 342370 399144 349838 399242
rect 350006 399144 357566 399242
rect 357734 399144 365202 399242
rect 365370 399144 372930 399242
rect 373098 399144 380658 399242
rect 380826 399144 388294 399242
rect 388462 399144 396022 399242
rect 396190 399144 398248 399242
rect 1398 856 398248 399144
rect 1398 800 2722 856
rect 2890 800 8334 856
rect 8502 800 13946 856
rect 14114 800 19558 856
rect 19726 800 25170 856
rect 25338 800 30874 856
rect 31042 800 36486 856
rect 36654 800 42098 856
rect 42266 800 47710 856
rect 47878 800 53414 856
rect 53582 800 59026 856
rect 59194 800 64638 856
rect 64806 800 70250 856
rect 70418 800 75954 856
rect 76122 800 81566 856
rect 81734 800 87178 856
rect 87346 800 92790 856
rect 92958 800 98494 856
rect 98662 800 104106 856
rect 104274 800 109718 856
rect 109886 800 115330 856
rect 115498 800 121034 856
rect 121202 800 126646 856
rect 126814 800 132258 856
rect 132426 800 137870 856
rect 138038 800 143482 856
rect 143650 800 149186 856
rect 149354 800 154798 856
rect 154966 800 160410 856
rect 160578 800 166022 856
rect 166190 800 171726 856
rect 171894 800 177338 856
rect 177506 800 182950 856
rect 183118 800 188562 856
rect 188730 800 194266 856
rect 194434 800 199878 856
rect 200046 800 205490 856
rect 205658 800 211102 856
rect 211270 800 216806 856
rect 216974 800 222418 856
rect 222586 800 228030 856
rect 228198 800 233642 856
rect 233810 800 239346 856
rect 239514 800 244958 856
rect 245126 800 250570 856
rect 250738 800 256182 856
rect 256350 800 261886 856
rect 262054 800 267498 856
rect 267666 800 273110 856
rect 273278 800 278722 856
rect 278890 800 284334 856
rect 284502 800 290038 856
rect 290206 800 295650 856
rect 295818 800 301262 856
rect 301430 800 306874 856
rect 307042 800 312578 856
rect 312746 800 318190 856
rect 318358 800 323802 856
rect 323970 800 329414 856
rect 329582 800 335118 856
rect 335286 800 340730 856
rect 340898 800 346342 856
rect 346510 800 351954 856
rect 352122 800 357658 856
rect 357826 800 363270 856
rect 363438 800 368882 856
rect 369050 800 374494 856
rect 374662 800 380198 856
rect 380366 800 385810 856
rect 385978 800 391422 856
rect 391590 800 397034 856
rect 397202 800 398248 856
<< metal3 >>
rect 0 396720 800 396840
rect 399200 396720 400000 396840
rect 0 390464 800 390584
rect 399200 390600 400000 390720
rect 399200 384480 400000 384600
rect 0 384208 800 384328
rect 399200 378360 400000 378480
rect 0 377952 800 378072
rect 399200 372104 400000 372224
rect 0 371696 800 371816
rect 399200 365984 400000 366104
rect 0 365440 800 365560
rect 399200 359864 400000 359984
rect 0 359184 800 359304
rect 399200 353744 400000 353864
rect 0 352928 800 353048
rect 399200 347488 400000 347608
rect 0 346672 800 346792
rect 399200 341368 400000 341488
rect 0 340416 800 340536
rect 399200 335248 400000 335368
rect 0 334160 800 334280
rect 399200 329128 400000 329248
rect 0 327904 800 328024
rect 399200 322872 400000 322992
rect 0 321648 800 321768
rect 399200 316752 400000 316872
rect 0 315392 800 315512
rect 399200 310632 400000 310752
rect 0 309136 800 309256
rect 399200 304512 400000 304632
rect 0 302880 800 303000
rect 399200 298256 400000 298376
rect 0 296624 800 296744
rect 399200 292136 400000 292256
rect 0 290368 800 290488
rect 399200 286016 400000 286136
rect 0 284112 800 284232
rect 399200 279896 400000 280016
rect 0 277856 800 277976
rect 399200 273640 400000 273760
rect 0 271600 800 271720
rect 399200 267520 400000 267640
rect 0 265480 800 265600
rect 399200 261400 400000 261520
rect 0 259224 800 259344
rect 399200 255280 400000 255400
rect 0 252968 800 253088
rect 399200 249024 400000 249144
rect 0 246712 800 246832
rect 399200 242904 400000 243024
rect 0 240456 800 240576
rect 399200 236784 400000 236904
rect 0 234200 800 234320
rect 399200 230664 400000 230784
rect 0 227944 800 228064
rect 399200 224408 400000 224528
rect 0 221688 800 221808
rect 399200 218288 400000 218408
rect 0 215432 800 215552
rect 399200 212168 400000 212288
rect 0 209176 800 209296
rect 399200 206048 400000 206168
rect 0 202920 800 203040
rect 399200 199792 400000 199912
rect 0 196664 800 196784
rect 399200 193672 400000 193792
rect 0 190408 800 190528
rect 399200 187552 400000 187672
rect 0 184152 800 184272
rect 399200 181432 400000 181552
rect 0 177896 800 178016
rect 399200 175176 400000 175296
rect 0 171640 800 171760
rect 399200 169056 400000 169176
rect 0 165384 800 165504
rect 399200 162936 400000 163056
rect 0 159128 800 159248
rect 399200 156816 400000 156936
rect 0 152872 800 152992
rect 399200 150560 400000 150680
rect 0 146616 800 146736
rect 399200 144440 400000 144560
rect 0 140360 800 140480
rect 399200 138320 400000 138440
rect 0 134240 800 134360
rect 399200 132200 400000 132320
rect 0 127984 800 128104
rect 399200 125944 400000 126064
rect 0 121728 800 121848
rect 399200 119824 400000 119944
rect 0 115472 800 115592
rect 399200 113704 400000 113824
rect 0 109216 800 109336
rect 399200 107584 400000 107704
rect 0 102960 800 103080
rect 399200 101328 400000 101448
rect 0 96704 800 96824
rect 399200 95208 400000 95328
rect 0 90448 800 90568
rect 399200 89088 400000 89208
rect 0 84192 800 84312
rect 399200 82968 400000 83088
rect 0 77936 800 78056
rect 399200 76712 400000 76832
rect 0 71680 800 71800
rect 399200 70592 400000 70712
rect 0 65424 800 65544
rect 399200 64472 400000 64592
rect 0 59168 800 59288
rect 399200 58352 400000 58472
rect 0 52912 800 53032
rect 399200 52096 400000 52216
rect 0 46656 800 46776
rect 399200 45976 400000 46096
rect 0 40400 800 40520
rect 399200 39856 400000 39976
rect 0 34144 800 34264
rect 399200 33736 400000 33856
rect 0 27888 800 28008
rect 399200 27480 400000 27600
rect 0 21632 800 21752
rect 399200 21360 400000 21480
rect 0 15376 800 15496
rect 399200 15240 400000 15360
rect 0 9120 800 9240
rect 399200 9120 400000 9240
rect 0 3000 800 3120
rect 399200 3000 400000 3120
<< obsm3 >>
rect 800 396920 399200 397697
rect 880 396640 399120 396920
rect 800 390800 399200 396640
rect 800 390664 399120 390800
rect 880 390520 399120 390664
rect 880 390384 399200 390520
rect 800 384680 399200 390384
rect 800 384408 399120 384680
rect 880 384400 399120 384408
rect 880 384128 399200 384400
rect 800 378560 399200 384128
rect 800 378280 399120 378560
rect 800 378152 399200 378280
rect 880 377872 399200 378152
rect 800 372304 399200 377872
rect 800 372024 399120 372304
rect 800 371896 399200 372024
rect 880 371616 399200 371896
rect 800 366184 399200 371616
rect 800 365904 399120 366184
rect 800 365640 399200 365904
rect 880 365360 399200 365640
rect 800 360064 399200 365360
rect 800 359784 399120 360064
rect 800 359384 399200 359784
rect 880 359104 399200 359384
rect 800 353944 399200 359104
rect 800 353664 399120 353944
rect 800 353128 399200 353664
rect 880 352848 399200 353128
rect 800 347688 399200 352848
rect 800 347408 399120 347688
rect 800 346872 399200 347408
rect 880 346592 399200 346872
rect 800 341568 399200 346592
rect 800 341288 399120 341568
rect 800 340616 399200 341288
rect 880 340336 399200 340616
rect 800 335448 399200 340336
rect 800 335168 399120 335448
rect 800 334360 399200 335168
rect 880 334080 399200 334360
rect 800 329328 399200 334080
rect 800 329048 399120 329328
rect 800 328104 399200 329048
rect 880 327824 399200 328104
rect 800 323072 399200 327824
rect 800 322792 399120 323072
rect 800 321848 399200 322792
rect 880 321568 399200 321848
rect 800 316952 399200 321568
rect 800 316672 399120 316952
rect 800 315592 399200 316672
rect 880 315312 399200 315592
rect 800 310832 399200 315312
rect 800 310552 399120 310832
rect 800 309336 399200 310552
rect 880 309056 399200 309336
rect 800 304712 399200 309056
rect 800 304432 399120 304712
rect 800 303080 399200 304432
rect 880 302800 399200 303080
rect 800 298456 399200 302800
rect 800 298176 399120 298456
rect 800 296824 399200 298176
rect 880 296544 399200 296824
rect 800 292336 399200 296544
rect 800 292056 399120 292336
rect 800 290568 399200 292056
rect 880 290288 399200 290568
rect 800 286216 399200 290288
rect 800 285936 399120 286216
rect 800 284312 399200 285936
rect 880 284032 399200 284312
rect 800 280096 399200 284032
rect 800 279816 399120 280096
rect 800 278056 399200 279816
rect 880 277776 399200 278056
rect 800 273840 399200 277776
rect 800 273560 399120 273840
rect 800 271800 399200 273560
rect 880 271520 399200 271800
rect 800 267720 399200 271520
rect 800 267440 399120 267720
rect 800 265680 399200 267440
rect 880 265400 399200 265680
rect 800 261600 399200 265400
rect 800 261320 399120 261600
rect 800 259424 399200 261320
rect 880 259144 399200 259424
rect 800 255480 399200 259144
rect 800 255200 399120 255480
rect 800 253168 399200 255200
rect 880 252888 399200 253168
rect 800 249224 399200 252888
rect 800 248944 399120 249224
rect 800 246912 399200 248944
rect 880 246632 399200 246912
rect 800 243104 399200 246632
rect 800 242824 399120 243104
rect 800 240656 399200 242824
rect 880 240376 399200 240656
rect 800 236984 399200 240376
rect 800 236704 399120 236984
rect 800 234400 399200 236704
rect 880 234120 399200 234400
rect 800 230864 399200 234120
rect 800 230584 399120 230864
rect 800 228144 399200 230584
rect 880 227864 399200 228144
rect 800 224608 399200 227864
rect 800 224328 399120 224608
rect 800 221888 399200 224328
rect 880 221608 399200 221888
rect 800 218488 399200 221608
rect 800 218208 399120 218488
rect 800 215632 399200 218208
rect 880 215352 399200 215632
rect 800 212368 399200 215352
rect 800 212088 399120 212368
rect 800 209376 399200 212088
rect 880 209096 399200 209376
rect 800 206248 399200 209096
rect 800 205968 399120 206248
rect 800 203120 399200 205968
rect 880 202840 399200 203120
rect 800 199992 399200 202840
rect 800 199712 399120 199992
rect 800 196864 399200 199712
rect 880 196584 399200 196864
rect 800 193872 399200 196584
rect 800 193592 399120 193872
rect 800 190608 399200 193592
rect 880 190328 399200 190608
rect 800 187752 399200 190328
rect 800 187472 399120 187752
rect 800 184352 399200 187472
rect 880 184072 399200 184352
rect 800 181632 399200 184072
rect 800 181352 399120 181632
rect 800 178096 399200 181352
rect 880 177816 399200 178096
rect 800 175376 399200 177816
rect 800 175096 399120 175376
rect 800 171840 399200 175096
rect 880 171560 399200 171840
rect 800 169256 399200 171560
rect 800 168976 399120 169256
rect 800 165584 399200 168976
rect 880 165304 399200 165584
rect 800 163136 399200 165304
rect 800 162856 399120 163136
rect 800 159328 399200 162856
rect 880 159048 399200 159328
rect 800 157016 399200 159048
rect 800 156736 399120 157016
rect 800 153072 399200 156736
rect 880 152792 399200 153072
rect 800 150760 399200 152792
rect 800 150480 399120 150760
rect 800 146816 399200 150480
rect 880 146536 399200 146816
rect 800 144640 399200 146536
rect 800 144360 399120 144640
rect 800 140560 399200 144360
rect 880 140280 399200 140560
rect 800 138520 399200 140280
rect 800 138240 399120 138520
rect 800 134440 399200 138240
rect 880 134160 399200 134440
rect 800 132400 399200 134160
rect 800 132120 399120 132400
rect 800 128184 399200 132120
rect 880 127904 399200 128184
rect 800 126144 399200 127904
rect 800 125864 399120 126144
rect 800 121928 399200 125864
rect 880 121648 399200 121928
rect 800 120024 399200 121648
rect 800 119744 399120 120024
rect 800 115672 399200 119744
rect 880 115392 399200 115672
rect 800 113904 399200 115392
rect 800 113624 399120 113904
rect 800 109416 399200 113624
rect 880 109136 399200 109416
rect 800 107784 399200 109136
rect 800 107504 399120 107784
rect 800 103160 399200 107504
rect 880 102880 399200 103160
rect 800 101528 399200 102880
rect 800 101248 399120 101528
rect 800 96904 399200 101248
rect 880 96624 399200 96904
rect 800 95408 399200 96624
rect 800 95128 399120 95408
rect 800 90648 399200 95128
rect 880 90368 399200 90648
rect 800 89288 399200 90368
rect 800 89008 399120 89288
rect 800 84392 399200 89008
rect 880 84112 399200 84392
rect 800 83168 399200 84112
rect 800 82888 399120 83168
rect 800 78136 399200 82888
rect 880 77856 399200 78136
rect 800 76912 399200 77856
rect 800 76632 399120 76912
rect 800 71880 399200 76632
rect 880 71600 399200 71880
rect 800 70792 399200 71600
rect 800 70512 399120 70792
rect 800 65624 399200 70512
rect 880 65344 399200 65624
rect 800 64672 399200 65344
rect 800 64392 399120 64672
rect 800 59368 399200 64392
rect 880 59088 399200 59368
rect 800 58552 399200 59088
rect 800 58272 399120 58552
rect 800 53112 399200 58272
rect 880 52832 399200 53112
rect 800 52296 399200 52832
rect 800 52016 399120 52296
rect 800 46856 399200 52016
rect 880 46576 399200 46856
rect 800 46176 399200 46576
rect 800 45896 399120 46176
rect 800 40600 399200 45896
rect 880 40320 399200 40600
rect 800 40056 399200 40320
rect 800 39776 399120 40056
rect 800 34344 399200 39776
rect 880 34064 399200 34344
rect 800 33936 399200 34064
rect 800 33656 399120 33936
rect 800 28088 399200 33656
rect 880 27808 399200 28088
rect 800 27680 399200 27808
rect 800 27400 399120 27680
rect 800 21832 399200 27400
rect 880 21560 399200 21832
rect 880 21552 399120 21560
rect 800 21280 399120 21552
rect 800 15576 399200 21280
rect 880 15440 399200 15576
rect 880 15296 399120 15440
rect 800 15160 399120 15296
rect 800 9320 399200 15160
rect 880 9040 399120 9320
rect 800 3200 399200 9040
rect 880 2920 399120 3200
rect 800 2143 399200 2920
<< metal4 >>
rect 4208 2128 4528 397712
rect 19568 2128 19888 397712
rect 34928 2128 35248 397712
rect 50288 2128 50608 397712
rect 65648 2128 65968 397712
rect 81008 2128 81328 397712
rect 96368 2128 96688 397712
rect 111728 2128 112048 397712
rect 127088 2128 127408 397712
rect 142448 2128 142768 397712
rect 157808 2128 158128 397712
rect 173168 2128 173488 397712
rect 188528 2128 188848 397712
rect 203888 2128 204208 397712
rect 219248 2128 219568 397712
rect 234608 2128 234928 397712
rect 249968 2128 250288 397712
rect 265328 2128 265648 397712
rect 280688 2128 281008 397712
rect 296048 2128 296368 397712
rect 311408 2128 311728 397712
rect 326768 2128 327088 397712
rect 342128 2128 342448 397712
rect 357488 2128 357808 397712
rect 372848 2128 373168 397712
rect 388208 2128 388528 397712
<< labels >>
rlabel metal2 s 3790 399200 3846 400000 6 clk
port 1 nsew signal input
rlabel metal3 s 399200 3000 400000 3120 6 external_interrupt
port 2 nsew signal input
rlabel metal3 s 399200 9120 400000 9240 6 l15_transducer_ack
port 3 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 l15_transducer_data_0[0]
port 4 nsew signal input
rlabel metal3 s 399200 70592 400000 70712 6 l15_transducer_data_0[10]
port 5 nsew signal input
rlabel metal2 s 119158 399200 119214 400000 6 l15_transducer_data_0[11]
port 6 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 l15_transducer_data_0[12]
port 7 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 l15_transducer_data_0[13]
port 8 nsew signal input
rlabel metal3 s 0 134240 800 134360 6 l15_transducer_data_0[14]
port 9 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 l15_transducer_data_0[15]
port 10 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 l15_transducer_data_0[16]
port 11 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 l15_transducer_data_0[17]
port 12 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 l15_transducer_data_0[18]
port 13 nsew signal input
rlabel metal3 s 0 177896 800 178016 6 l15_transducer_data_0[19]
port 14 nsew signal input
rlabel metal3 s 399200 21360 400000 21480 6 l15_transducer_data_0[1]
port 15 nsew signal input
rlabel metal3 s 399200 150560 400000 150680 6 l15_transducer_data_0[20]
port 16 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 l15_transducer_data_0[21]
port 17 nsew signal input
rlabel metal3 s 0 202920 800 203040 6 l15_transducer_data_0[22]
port 18 nsew signal input
rlabel metal3 s 0 215432 800 215552 6 l15_transducer_data_0[23]
port 19 nsew signal input
rlabel metal3 s 0 227944 800 228064 6 l15_transducer_data_0[24]
port 20 nsew signal input
rlabel metal3 s 0 240456 800 240576 6 l15_transducer_data_0[25]
port 21 nsew signal input
rlabel metal3 s 399200 199792 400000 199912 6 l15_transducer_data_0[26]
port 22 nsew signal input
rlabel metal3 s 399200 212168 400000 212288 6 l15_transducer_data_0[27]
port 23 nsew signal input
rlabel metal2 s 180706 399200 180762 400000 6 l15_transducer_data_0[28]
port 24 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 l15_transducer_data_0[29]
port 25 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 l15_transducer_data_0[2]
port 26 nsew signal input
rlabel metal2 s 203798 399200 203854 400000 6 l15_transducer_data_0[30]
port 27 nsew signal input
rlabel metal2 s 211158 0 211214 800 6 l15_transducer_data_0[31]
port 28 nsew signal input
rlabel metal3 s 0 265480 800 265600 6 l15_transducer_data_0[32]
port 29 nsew signal input
rlabel metal3 s 399200 249024 400000 249144 6 l15_transducer_data_0[33]
port 30 nsew signal input
rlabel metal3 s 0 277856 800 277976 6 l15_transducer_data_0[34]
port 31 nsew signal input
rlabel metal3 s 0 284112 800 284232 6 l15_transducer_data_0[35]
port 32 nsew signal input
rlabel metal3 s 399200 261400 400000 261520 6 l15_transducer_data_0[36]
port 33 nsew signal input
rlabel metal3 s 0 315392 800 315512 6 l15_transducer_data_0[37]
port 34 nsew signal input
rlabel metal3 s 399200 286016 400000 286136 6 l15_transducer_data_0[38]
port 35 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 l15_transducer_data_0[39]
port 36 nsew signal input
rlabel metal2 s 49882 399200 49938 400000 6 l15_transducer_data_0[3]
port 37 nsew signal input
rlabel metal3 s 399200 298256 400000 298376 6 l15_transducer_data_0[40]
port 38 nsew signal input
rlabel metal3 s 0 340416 800 340536 6 l15_transducer_data_0[41]
port 39 nsew signal input
rlabel metal2 s 261942 0 261998 800 6 l15_transducer_data_0[42]
port 40 nsew signal input
rlabel metal3 s 399200 310632 400000 310752 6 l15_transducer_data_0[43]
port 41 nsew signal input
rlabel metal2 s 278778 0 278834 800 6 l15_transducer_data_0[44]
port 42 nsew signal input
rlabel metal3 s 0 352928 800 353048 6 l15_transducer_data_0[45]
port 43 nsew signal input
rlabel metal2 s 284390 0 284446 800 6 l15_transducer_data_0[46]
port 44 nsew signal input
rlabel metal2 s 290094 0 290150 800 6 l15_transducer_data_0[47]
port 45 nsew signal input
rlabel metal2 s 296074 399200 296130 400000 6 l15_transducer_data_0[48]
port 46 nsew signal input
rlabel metal2 s 303802 399200 303858 400000 6 l15_transducer_data_0[49]
port 47 nsew signal input
rlabel metal2 s 72974 399200 73030 400000 6 l15_transducer_data_0[4]
port 48 nsew signal input
rlabel metal2 s 312634 0 312690 800 6 l15_transducer_data_0[50]
port 49 nsew signal input
rlabel metal2 s 318246 0 318302 800 6 l15_transducer_data_0[51]
port 50 nsew signal input
rlabel metal2 s 342258 399200 342314 400000 6 l15_transducer_data_0[52]
port 51 nsew signal input
rlabel metal2 s 323858 0 323914 800 6 l15_transducer_data_0[53]
port 52 nsew signal input
rlabel metal3 s 0 377952 800 378072 6 l15_transducer_data_0[54]
port 53 nsew signal input
rlabel metal2 s 340786 0 340842 800 6 l15_transducer_data_0[55]
port 54 nsew signal input
rlabel metal2 s 352010 0 352066 800 6 l15_transducer_data_0[56]
port 55 nsew signal input
rlabel metal2 s 363326 0 363382 800 6 l15_transducer_data_0[57]
port 56 nsew signal input
rlabel metal3 s 399200 365984 400000 366104 6 l15_transducer_data_0[58]
port 57 nsew signal input
rlabel metal2 s 365258 399200 365314 400000 6 l15_transducer_data_0[59]
port 58 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 l15_transducer_data_0[5]
port 59 nsew signal input
rlabel metal2 s 388350 399200 388406 400000 6 l15_transducer_data_0[60]
port 60 nsew signal input
rlabel metal2 s 380254 0 380310 800 6 l15_transducer_data_0[61]
port 61 nsew signal input
rlabel metal3 s 399200 372104 400000 372224 6 l15_transducer_data_0[62]
port 62 nsew signal input
rlabel metal2 s 397090 0 397146 800 6 l15_transducer_data_0[63]
port 63 nsew signal input
rlabel metal2 s 88338 399200 88394 400000 6 l15_transducer_data_0[6]
port 64 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 l15_transducer_data_0[7]
port 65 nsew signal input
rlabel metal2 s 96066 399200 96122 400000 6 l15_transducer_data_0[8]
port 66 nsew signal input
rlabel metal2 s 103794 399200 103850 400000 6 l15_transducer_data_0[9]
port 67 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 l15_transducer_data_1[0]
port 68 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 l15_transducer_data_1[10]
port 69 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 l15_transducer_data_1[11]
port 70 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 l15_transducer_data_1[12]
port 71 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 l15_transducer_data_1[13]
port 72 nsew signal input
rlabel metal3 s 399200 101328 400000 101448 6 l15_transducer_data_1[14]
port 73 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 l15_transducer_data_1[15]
port 74 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 l15_transducer_data_1[16]
port 75 nsew signal input
rlabel metal2 s 126794 399200 126850 400000 6 l15_transducer_data_1[17]
port 76 nsew signal input
rlabel metal2 s 142250 399200 142306 400000 6 l15_transducer_data_1[18]
port 77 nsew signal input
rlabel metal3 s 399200 138320 400000 138440 6 l15_transducer_data_1[19]
port 78 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 l15_transducer_data_1[1]
port 79 nsew signal input
rlabel metal3 s 0 184152 800 184272 6 l15_transducer_data_1[20]
port 80 nsew signal input
rlabel metal3 s 399200 169056 400000 169176 6 l15_transducer_data_1[21]
port 81 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 l15_transducer_data_1[22]
port 82 nsew signal input
rlabel metal3 s 0 221688 800 221808 6 l15_transducer_data_1[23]
port 83 nsew signal input
rlabel metal3 s 0 234200 800 234320 6 l15_transducer_data_1[24]
port 84 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 l15_transducer_data_1[25]
port 85 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 l15_transducer_data_1[26]
port 86 nsew signal input
rlabel metal2 s 172978 399200 173034 400000 6 l15_transducer_data_1[27]
port 87 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 l15_transducer_data_1[28]
port 88 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 l15_transducer_data_1[29]
port 89 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 l15_transducer_data_1[2]
port 90 nsew signal input
rlabel metal2 s 211434 399200 211490 400000 6 l15_transducer_data_1[30]
port 91 nsew signal input
rlabel metal3 s 0 259224 800 259344 6 l15_transducer_data_1[31]
port 92 nsew signal input
rlabel metal3 s 0 271600 800 271720 6 l15_transducer_data_1[32]
port 93 nsew signal input
rlabel metal2 s 226798 399200 226854 400000 6 l15_transducer_data_1[33]
port 94 nsew signal input
rlabel metal2 s 234526 399200 234582 400000 6 l15_transducer_data_1[34]
port 95 nsew signal input
rlabel metal3 s 0 290368 800 290488 6 l15_transducer_data_1[35]
port 96 nsew signal input
rlabel metal3 s 0 302880 800 303000 6 l15_transducer_data_1[36]
port 97 nsew signal input
rlabel metal3 s 399200 273640 400000 273760 6 l15_transducer_data_1[37]
port 98 nsew signal input
rlabel metal3 s 399200 292136 400000 292256 6 l15_transducer_data_1[38]
port 99 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 l15_transducer_data_1[39]
port 100 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 l15_transducer_data_1[3]
port 101 nsew signal input
rlabel metal3 s 0 334160 800 334280 6 l15_transducer_data_1[40]
port 102 nsew signal input
rlabel metal3 s 399200 304512 400000 304632 6 l15_transducer_data_1[41]
port 103 nsew signal input
rlabel metal2 s 267554 0 267610 800 6 l15_transducer_data_1[42]
port 104 nsew signal input
rlabel metal3 s 0 346672 800 346792 6 l15_transducer_data_1[43]
port 105 nsew signal input
rlabel metal2 s 272982 399200 273038 400000 6 l15_transducer_data_1[44]
port 106 nsew signal input
rlabel metal3 s 0 359184 800 359304 6 l15_transducer_data_1[45]
port 107 nsew signal input
rlabel metal3 s 0 365440 800 365560 6 l15_transducer_data_1[46]
port 108 nsew signal input
rlabel metal2 s 295706 0 295762 800 6 l15_transducer_data_1[47]
port 109 nsew signal input
rlabel metal2 s 301318 0 301374 800 6 l15_transducer_data_1[48]
port 110 nsew signal input
rlabel metal2 s 311438 399200 311494 400000 6 l15_transducer_data_1[49]
port 111 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 l15_transducer_data_1[4]
port 112 nsew signal input
rlabel metal2 s 319166 399200 319222 400000 6 l15_transducer_data_1[50]
port 113 nsew signal input
rlabel metal2 s 334530 399200 334586 400000 6 l15_transducer_data_1[51]
port 114 nsew signal input
rlabel metal3 s 399200 347488 400000 347608 6 l15_transducer_data_1[52]
port 115 nsew signal input
rlabel metal2 s 329470 0 329526 800 6 l15_transducer_data_1[53]
port 116 nsew signal input
rlabel metal2 s 349894 399200 349950 400000 6 l15_transducer_data_1[54]
port 117 nsew signal input
rlabel metal2 s 357622 399200 357678 400000 6 l15_transducer_data_1[55]
port 118 nsew signal input
rlabel metal3 s 399200 353744 400000 353864 6 l15_transducer_data_1[56]
port 119 nsew signal input
rlabel metal3 s 399200 359864 400000 359984 6 l15_transducer_data_1[57]
port 120 nsew signal input
rlabel metal2 s 374550 0 374606 800 6 l15_transducer_data_1[58]
port 121 nsew signal input
rlabel metal2 s 372986 399200 373042 400000 6 l15_transducer_data_1[59]
port 122 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 l15_transducer_data_1[5]
port 123 nsew signal input
rlabel metal2 s 396078 399200 396134 400000 6 l15_transducer_data_1[60]
port 124 nsew signal input
rlabel metal2 s 385866 0 385922 800 6 l15_transducer_data_1[61]
port 125 nsew signal input
rlabel metal3 s 399200 378360 400000 378480 6 l15_transducer_data_1[62]
port 126 nsew signal input
rlabel metal3 s 399200 390600 400000 390720 6 l15_transducer_data_1[63]
port 127 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 l15_transducer_data_1[6]
port 128 nsew signal input
rlabel metal3 s 0 96704 800 96824 6 l15_transducer_data_1[7]
port 129 nsew signal input
rlabel metal3 s 399200 45976 400000 46096 6 l15_transducer_data_1[8]
port 130 nsew signal input
rlabel metal3 s 399200 52096 400000 52216 6 l15_transducer_data_1[9]
port 131 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 l15_transducer_header_ack
port 132 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 l15_transducer_returntype[0]
port 133 nsew signal input
rlabel metal3 s 399200 27480 400000 27600 6 l15_transducer_returntype[1]
port 134 nsew signal input
rlabel metal2 s 34518 399200 34574 400000 6 l15_transducer_returntype[2]
port 135 nsew signal input
rlabel metal2 s 57610 399200 57666 400000 6 l15_transducer_returntype[3]
port 136 nsew signal input
rlabel metal2 s 11426 399200 11482 400000 6 l15_transducer_val
port 137 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 nrst
port 138 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 transducer_l15_address[0]
port 139 nsew signal output
rlabel metal2 s 111430 399200 111486 400000 6 transducer_l15_address[10]
port 140 nsew signal output
rlabel metal3 s 399200 76712 400000 76832 6 transducer_l15_address[11]
port 141 nsew signal output
rlabel metal3 s 399200 89088 400000 89208 6 transducer_l15_address[12]
port 142 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 transducer_l15_address[13]
port 143 nsew signal output
rlabel metal3 s 399200 107584 400000 107704 6 transducer_l15_address[14]
port 144 nsew signal output
rlabel metal3 s 399200 113704 400000 113824 6 transducer_l15_address[15]
port 145 nsew signal output
rlabel metal3 s 399200 125944 400000 126064 6 transducer_l15_address[16]
port 146 nsew signal output
rlabel metal3 s 0 165384 800 165504 6 transducer_l15_address[17]
port 147 nsew signal output
rlabel metal3 s 399200 132200 400000 132320 6 transducer_l15_address[18]
port 148 nsew signal output
rlabel metal3 s 399200 144440 400000 144560 6 transducer_l15_address[19]
port 149 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 transducer_l15_address[1]
port 150 nsew signal output
rlabel metal3 s 399200 156816 400000 156936 6 transducer_l15_address[20]
port 151 nsew signal output
rlabel metal3 s 399200 175176 400000 175296 6 transducer_l15_address[21]
port 152 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 transducer_l15_address[22]
port 153 nsew signal output
rlabel metal2 s 157614 399200 157670 400000 6 transducer_l15_address[23]
port 154 nsew signal output
rlabel metal3 s 399200 187552 400000 187672 6 transducer_l15_address[24]
port 155 nsew signal output
rlabel metal3 s 399200 193672 400000 193792 6 transducer_l15_address[25]
port 156 nsew signal output
rlabel metal3 s 0 246712 800 246832 6 transducer_l15_address[26]
port 157 nsew signal output
rlabel metal3 s 399200 218288 400000 218408 6 transducer_l15_address[27]
port 158 nsew signal output
rlabel metal3 s 399200 224408 400000 224528 6 transducer_l15_address[28]
port 159 nsew signal output
rlabel metal2 s 188342 399200 188398 400000 6 transducer_l15_address[29]
port 160 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 transducer_l15_address[2]
port 161 nsew signal output
rlabel metal2 s 205546 0 205602 800 6 transducer_l15_address[30]
port 162 nsew signal output
rlabel metal3 s 399200 236784 400000 236904 6 transducer_l15_address[31]
port 163 nsew signal output
rlabel metal2 s 216862 0 216918 800 6 transducer_l15_address[32]
port 164 nsew signal output
rlabel metal3 s 399200 255280 400000 255400 6 transducer_l15_address[33]
port 165 nsew signal output
rlabel metal2 s 228086 0 228142 800 6 transducer_l15_address[34]
port 166 nsew signal output
rlabel metal3 s 0 296624 800 296744 6 transducer_l15_address[35]
port 167 nsew signal output
rlabel metal3 s 399200 267520 400000 267640 6 transducer_l15_address[36]
port 168 nsew signal output
rlabel metal3 s 399200 279896 400000 280016 6 transducer_l15_address[37]
port 169 nsew signal output
rlabel metal2 s 233698 0 233754 800 6 transducer_l15_address[38]
port 170 nsew signal output
rlabel metal3 s 0 327904 800 328024 6 transducer_l15_address[39]
port 171 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 transducer_l15_address[3]
port 172 nsew signal output
rlabel metal2 s 80702 399200 80758 400000 6 transducer_l15_address[4]
port 173 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 transducer_l15_address[5]
port 174 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 transducer_l15_address[6]
port 175 nsew signal output
rlabel metal3 s 0 102960 800 103080 6 transducer_l15_address[7]
port 176 nsew signal output
rlabel metal3 s 0 109216 800 109336 6 transducer_l15_address[8]
port 177 nsew signal output
rlabel metal3 s 399200 58352 400000 58472 6 transducer_l15_address[9]
port 178 nsew signal output
rlabel metal2 s 19154 399200 19210 400000 6 transducer_l15_data[0]
port 179 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 transducer_l15_data[10]
port 180 nsew signal output
rlabel metal3 s 399200 82968 400000 83088 6 transducer_l15_data[11]
port 181 nsew signal output
rlabel metal3 s 399200 95208 400000 95328 6 transducer_l15_data[12]
port 182 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 transducer_l15_data[13]
port 183 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 transducer_l15_data[14]
port 184 nsew signal output
rlabel metal3 s 399200 119824 400000 119944 6 transducer_l15_data[15]
port 185 nsew signal output
rlabel metal3 s 0 152872 800 152992 6 transducer_l15_data[16]
port 186 nsew signal output
rlabel metal2 s 134522 399200 134578 400000 6 transducer_l15_data[17]
port 187 nsew signal output
rlabel metal3 s 0 171640 800 171760 6 transducer_l15_data[18]
port 188 nsew signal output
rlabel metal2 s 149886 399200 149942 400000 6 transducer_l15_data[19]
port 189 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 transducer_l15_data[1]
port 190 nsew signal output
rlabel metal3 s 399200 162936 400000 163056 6 transducer_l15_data[20]
port 191 nsew signal output
rlabel metal3 s 0 196664 800 196784 6 transducer_l15_data[21]
port 192 nsew signal output
rlabel metal3 s 0 209176 800 209296 6 transducer_l15_data[22]
port 193 nsew signal output
rlabel metal3 s 399200 181432 400000 181552 6 transducer_l15_data[23]
port 194 nsew signal output
rlabel metal2 s 165250 399200 165306 400000 6 transducer_l15_data[24]
port 195 nsew signal output
rlabel metal2 s 171782 0 171838 800 6 transducer_l15_data[25]
port 196 nsew signal output
rlabel metal3 s 399200 206048 400000 206168 6 transducer_l15_data[26]
port 197 nsew signal output
rlabel metal2 s 183006 0 183062 800 6 transducer_l15_data[27]
port 198 nsew signal output
rlabel metal3 s 399200 230664 400000 230784 6 transducer_l15_data[28]
port 199 nsew signal output
rlabel metal2 s 196070 399200 196126 400000 6 transducer_l15_data[29]
port 200 nsew signal output
rlabel metal2 s 42246 399200 42302 400000 6 transducer_l15_data[2]
port 201 nsew signal output
rlabel metal3 s 0 252968 800 253088 6 transducer_l15_data[30]
port 202 nsew signal output
rlabel metal2 s 219162 399200 219218 400000 6 transducer_l15_data[31]
port 203 nsew signal output
rlabel metal3 s 399200 242904 400000 243024 6 transducer_l15_data[32]
port 204 nsew signal output
rlabel metal2 s 222474 0 222530 800 6 transducer_l15_data[33]
port 205 nsew signal output
rlabel metal2 s 242254 399200 242310 400000 6 transducer_l15_data[34]
port 206 nsew signal output
rlabel metal2 s 249890 399200 249946 400000 6 transducer_l15_data[35]
port 207 nsew signal output
rlabel metal3 s 0 309136 800 309256 6 transducer_l15_data[36]
port 208 nsew signal output
rlabel metal3 s 0 321648 800 321768 6 transducer_l15_data[37]
port 209 nsew signal output
rlabel metal2 s 239402 0 239458 800 6 transducer_l15_data[38]
port 210 nsew signal output
rlabel metal2 s 256238 0 256294 800 6 transducer_l15_data[39]
port 211 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 transducer_l15_data[3]
port 212 nsew signal output
rlabel metal2 s 257618 399200 257674 400000 6 transducer_l15_data[40]
port 213 nsew signal output
rlabel metal2 s 265254 399200 265310 400000 6 transducer_l15_data[41]
port 214 nsew signal output
rlabel metal2 s 273166 0 273222 800 6 transducer_l15_data[42]
port 215 nsew signal output
rlabel metal3 s 399200 316752 400000 316872 6 transducer_l15_data[43]
port 216 nsew signal output
rlabel metal2 s 280710 399200 280766 400000 6 transducer_l15_data[44]
port 217 nsew signal output
rlabel metal3 s 399200 322872 400000 322992 6 transducer_l15_data[45]
port 218 nsew signal output
rlabel metal3 s 399200 329128 400000 329248 6 transducer_l15_data[46]
port 219 nsew signal output
rlabel metal2 s 288346 399200 288402 400000 6 transducer_l15_data[47]
port 220 nsew signal output
rlabel metal3 s 399200 335248 400000 335368 6 transducer_l15_data[48]
port 221 nsew signal output
rlabel metal2 s 306930 0 306986 800 6 transducer_l15_data[49]
port 222 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 transducer_l15_data[4]
port 223 nsew signal output
rlabel metal2 s 326802 399200 326858 400000 6 transducer_l15_data[50]
port 224 nsew signal output
rlabel metal3 s 399200 341368 400000 341488 6 transducer_l15_data[51]
port 225 nsew signal output
rlabel metal3 s 0 371696 800 371816 6 transducer_l15_data[52]
port 226 nsew signal output
rlabel metal2 s 335174 0 335230 800 6 transducer_l15_data[53]
port 227 nsew signal output
rlabel metal3 s 0 384208 800 384328 6 transducer_l15_data[54]
port 228 nsew signal output
rlabel metal2 s 346398 0 346454 800 6 transducer_l15_data[55]
port 229 nsew signal output
rlabel metal2 s 357714 0 357770 800 6 transducer_l15_data[56]
port 230 nsew signal output
rlabel metal2 s 368938 0 368994 800 6 transducer_l15_data[57]
port 231 nsew signal output
rlabel metal3 s 0 390464 800 390584 6 transducer_l15_data[58]
port 232 nsew signal output
rlabel metal2 s 380714 399200 380770 400000 6 transducer_l15_data[59]
port 233 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 transducer_l15_data[5]
port 234 nsew signal output
rlabel metal3 s 0 396720 800 396840 6 transducer_l15_data[60]
port 235 nsew signal output
rlabel metal2 s 391478 0 391534 800 6 transducer_l15_data[61]
port 236 nsew signal output
rlabel metal3 s 399200 384480 400000 384600 6 transducer_l15_data[62]
port 237 nsew signal output
rlabel metal3 s 399200 396720 400000 396840 6 transducer_l15_data[63]
port 238 nsew signal output
rlabel metal3 s 0 84192 800 84312 6 transducer_l15_data[6]
port 239 nsew signal output
rlabel metal3 s 399200 39856 400000 39976 6 transducer_l15_data[7]
port 240 nsew signal output
rlabel metal3 s 0 115472 800 115592 6 transducer_l15_data[8]
port 241 nsew signal output
rlabel metal3 s 399200 64472 400000 64592 6 transducer_l15_data[9]
port 242 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 transducer_l15_req_ack
port 243 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 transducer_l15_rqtype[0]
port 244 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 transducer_l15_rqtype[1]
port 245 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 transducer_l15_rqtype[2]
port 246 nsew signal output
rlabel metal2 s 65246 399200 65302 400000 6 transducer_l15_rqtype[3]
port 247 nsew signal output
rlabel metal3 s 399200 33736 400000 33856 6 transducer_l15_rqtype[4]
port 248 nsew signal output
rlabel metal3 s 399200 15240 400000 15360 6 transducer_l15_size[0]
port 249 nsew signal output
rlabel metal2 s 26790 399200 26846 400000 6 transducer_l15_size[1]
port 250 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 transducer_l15_size[2]
port 251 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 transducer_l15_val
port 252 nsew signal output
rlabel metal4 s 4208 2128 4528 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 34928 2128 35248 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 65648 2128 65968 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 96368 2128 96688 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 127088 2128 127408 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 157808 2128 158128 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 188528 2128 188848 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 219248 2128 219568 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 249968 2128 250288 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 280688 2128 281008 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 311408 2128 311728 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 342128 2128 342448 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 372848 2128 373168 397712 6 vccd1
port 253 nsew power input
rlabel metal4 s 19568 2128 19888 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 50288 2128 50608 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 81008 2128 81328 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 111728 2128 112048 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 142448 2128 142768 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 173168 2128 173488 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 203888 2128 204208 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 234608 2128 234928 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 265328 2128 265648 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 296048 2128 296368 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 326768 2128 327088 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 357488 2128 357808 397712 6 vssd1
port 254 nsew ground input
rlabel metal4 s 388208 2128 388528 397712 6 vssd1
port 254 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 400000 400000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 43817766
string GDS_FILE /home/younis/caravel_tutorial/caravel_example/openlane/core/runs/core/results/finishing/core.magic.gds
string GDS_START 475516
<< end >>

